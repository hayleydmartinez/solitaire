module solitaire(clk, rst) begin
    // code here
endmodule